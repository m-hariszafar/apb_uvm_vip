interface apb_interface;
  logic pclk;
  logic presetn;
  logic [31:0] padder;
  logic pselx;
  logic penable;
  logic pwrite;
  logic [31:0] pwdata; 
  logic pready;
  logic [31:0] prdata;
  logic pslverr;

endinterface
