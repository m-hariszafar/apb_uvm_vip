package apb_package;

  import uvm_pkg::*;
    `include "tb/sequences/apb_transaction.sv"
	`include "tb/sequences/apb_sequences.sv"
    `include "tb/sequences/apb_wr_sequence.sv"
    `include "tb/sequences/apb_rd_sequence.sv"
    `include "tb/sequences/apb_sequencer.sv"
	`include "tb/agent/apb_driver.sv"
	`include "tb/agent/apb_coverage.sv"
	`include "tb/agent/apb_monitor.sv"
	`include "tb/agent/apb_agent.sv"
	`include "tb/env/apb_scoreboard.sv"
	`include "tb/env/apb_env.sv"
	`include "tb/test/apb_test.sv"
endpackage
